`define VLIB_BYPASS_POWER_CG
`define NV_FPGA_FIFOGEN
`define FIFOGEN_MASTER_CLK_GATING_DISABLED
`define FPGA
`define SYNTHESIS

// ================================================================
// NVDLA Open Source Project
//
// Copyright(c) 2016 - 2017 NVIDIA Corporation. Licensed under the
// NVDLA Open Hardware License; Check "LICENSE" which comes with
// this distribution for more information.
// ================================================================
// File Name: HLS_uint16_to_fp17.v
module UINT16_TO_FP17_mgc_in_wire_wait_v1 (ld, vd, d, lz, vz, z);
  parameter integer rscid = 1;
  parameter integer width = 8;
  input ld;
  output vd;
  output [width-1:0] d;
  output lz;
  input vz;
  input [width-1:0] z;
  wire vd;
  wire [width-1:0] d;
  wire lz;
  assign d = z;
  assign lz = ld;
  assign vd = vz;
endmodule
//------> /home/tools/calypto/catapult-10.0-264918/Mgc_home/pkgs/siflibs/UINT16_TO_FP17_mgc_out_stdreg_wait_v1.v
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
// All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------
module UINT16_TO_FP17_mgc_out_stdreg_wait_v1 (ld, vd, d, lz, vz, z);
  parameter integer rscid = 1;
  parameter integer width = 8;
  input ld;
  output vd;
  input [width-1:0] d;
  output lz;
  input vz;
  output [width-1:0] z;
  wire vd;
  wire lz;
  wire [width-1:0] z;
  assign z = d;
  assign lz = ld;
  assign vd = vz;
endmodule
//------> /home/tools/calypto/catapult-10.0-264918/Mgc_home/pkgs/siflibs/mgc_shift_l_beh_v4.v
module UINT16_TO_FP17_mgc_shift_l_v4(a,s,z);
   parameter width_a = 4;
   parameter signd_a = 1;
   parameter width_s = 2;
   parameter width_z = 8;
   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;
   generate
   if (signd_a)
   begin: SIGNED
      assign z = fshl_u(a,s,a[width_a-1]);
   end
   else
   begin: UNSIGNED
      assign z = fshl_u(a,s,1'b0);
   end
   endgenerate
//Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 = result[olen-1:0];
      end
   endfunction // fshl_u
//Shift-left - unsigned shift argument
   function [width_z-1:0] fshl_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      fshl_u = fshl_u_1({sbit,arg1} ,arg2, sbit);
   endfunction // fshl_u
endmodule
//------> ../td_ccore_solutions/leading_sign_16_0_584ce9c19228fa5400845cefe3e6770649bb_0/rtl.v
// ----------------------------------------------------------------------
// HLS HDL: Verilog Netlister
// HLS Version: 10.0/264918 Production Release
// HLS Date: Mon Aug 8 13:35:54 PDT 2016
//
// Generated by: ezhang@hk-sim-10-176
// Generated date: Wed Nov 23 14:25:06 2016
// ----------------------------------------------------------------------
//
// ------------------------------------------------------------------
// Design Unit: UINT16_TO_FP17_leading_sign_16_0
// ------------------------------------------------------------------
module UINT16_TO_FP17_leading_sign_16_0 (
  mantissa, rtn
);
  input [15:0] mantissa;
  output [4:0] rtn;
// Interconnect Declarations
  wire IntLeadZero_16U_leading_sign_16_0_rtn_wrs_c_6_2_sdt_2;
  wire IntLeadZero_16U_leading_sign_16_0_rtn_wrs_c_18_3_sdt_3;
  wire IntLeadZero_16U_leading_sign_16_0_rtn_wrs_c_26_2_sdt_2;
  wire IntLeadZero_16U_leading_sign_16_0_rtn_wrs_c_44_4_sdt_4;
  wire IntLeadZero_16U_leading_sign_16_0_rtn_wrs_c_6_2_sdt_1;
  wire IntLeadZero_16U_leading_sign_16_0_rtn_wrs_c_14_2_sdt_1;
  wire IntLeadZero_16U_leading_sign_16_0_rtn_wrs_c_26_2_sdt_1;
  wire IntLeadZero_16U_leading_sign_16_0_rtn_wrs_c_34_2_sdt_1;
  wire c_h_1_2;
  wire c_h_1_5;
  wire c_h_1_6;
  wire[3:0] IntLeadZero_16U_leading_sign_16_0_rtn_IntLeadZero_16U_leading_sign_16_0_rtn_and_nl;
  wire[0:0] IntLeadZero_16U_leading_sign_16_0_rtn_and_55_nl;
  wire[0:0] IntLeadZero_16U_leading_sign_16_0_rtn_and_53_nl;
  wire[0:0] IntLeadZero_16U_leading_sign_16_0_rtn_and_60_nl;
  wire[0:0] IntLeadZero_16U_leading_sign_16_0_rtn_not_nl;
// Interconnect Declarations for Component Instantiations
  assign IntLeadZero_16U_leading_sign_16_0_rtn_wrs_c_6_2_sdt_2 = ~((mantissa[13:12]!=2'b00));
  assign IntLeadZero_16U_leading_sign_16_0_rtn_wrs_c_6_2_sdt_1 = ~((mantissa[15:14]!=2'b00));
  assign IntLeadZero_16U_leading_sign_16_0_rtn_wrs_c_14_2_sdt_1 = ~((mantissa[11:10]!=2'b00));
  assign c_h_1_2 = IntLeadZero_16U_leading_sign_16_0_rtn_wrs_c_6_2_sdt_1 & IntLeadZero_16U_leading_sign_16_0_rtn_wrs_c_6_2_sdt_2;
  assign IntLeadZero_16U_leading_sign_16_0_rtn_wrs_c_18_3_sdt_3 = (mantissa[9:8]==2'b00)
      & IntLeadZero_16U_leading_sign_16_0_rtn_wrs_c_14_2_sdt_1;
  assign IntLeadZero_16U_leading_sign_16_0_rtn_wrs_c_26_2_sdt_2 = ~((mantissa[5:4]!=2'b00));
  assign IntLeadZero_16U_leading_sign_16_0_rtn_wrs_c_26_2_sdt_1 = ~((mantissa[7:6]!=2'b00));
  assign IntLeadZero_16U_leading_sign_16_0_rtn_wrs_c_34_2_sdt_1 = ~((mantissa[3:2]!=2'b00));
  assign c_h_1_5 = IntLeadZero_16U_leading_sign_16_0_rtn_wrs_c_26_2_sdt_1 & IntLeadZero_16U_leading_sign_16_0_rtn_wrs_c_26_2_sdt_2;
  assign c_h_1_6 = c_h_1_2 & IntLeadZero_16U_leading_sign_16_0_rtn_wrs_c_18_3_sdt_3;
  assign IntLeadZero_16U_leading_sign_16_0_rtn_wrs_c_44_4_sdt_4 = (mantissa[1:0]==2'b00)
      & IntLeadZero_16U_leading_sign_16_0_rtn_wrs_c_34_2_sdt_1 & c_h_1_5 & c_h_1_6;
  assign IntLeadZero_16U_leading_sign_16_0_rtn_and_55_nl = c_h_1_2 & (c_h_1_5 | (~
      IntLeadZero_16U_leading_sign_16_0_rtn_wrs_c_18_3_sdt_3));
  assign IntLeadZero_16U_leading_sign_16_0_rtn_and_53_nl = IntLeadZero_16U_leading_sign_16_0_rtn_wrs_c_6_2_sdt_1
      & (IntLeadZero_16U_leading_sign_16_0_rtn_wrs_c_14_2_sdt_1 | (~ IntLeadZero_16U_leading_sign_16_0_rtn_wrs_c_6_2_sdt_2))
      & (~((~(IntLeadZero_16U_leading_sign_16_0_rtn_wrs_c_26_2_sdt_1 & (IntLeadZero_16U_leading_sign_16_0_rtn_wrs_c_34_2_sdt_1
      | (~ IntLeadZero_16U_leading_sign_16_0_rtn_wrs_c_26_2_sdt_2)))) & c_h_1_6));
  assign IntLeadZero_16U_leading_sign_16_0_rtn_and_60_nl = (~((mantissa[15]) | (~((mantissa[14:13]!=2'b01)))))
      & (~(((mantissa[11]) | (~((mantissa[10:9]!=2'b01)))) & c_h_1_2)) & (~((~((~((mantissa[7])
      | (~((mantissa[6:5]!=2'b01))))) & (~(((mantissa[3]) | (~((mantissa[2:1]!=2'b01))))
      & c_h_1_5)))) & c_h_1_6));
  assign IntLeadZero_16U_leading_sign_16_0_rtn_not_nl = ~ IntLeadZero_16U_leading_sign_16_0_rtn_wrs_c_44_4_sdt_4;
  assign IntLeadZero_16U_leading_sign_16_0_rtn_IntLeadZero_16U_leading_sign_16_0_rtn_and_nl
      = MUX_v_4_2_2(4'b0000, ({c_h_1_6 , (IntLeadZero_16U_leading_sign_16_0_rtn_and_55_nl)
      , (IntLeadZero_16U_leading_sign_16_0_rtn_and_53_nl) , (IntLeadZero_16U_leading_sign_16_0_rtn_and_60_nl)}),
      (IntLeadZero_16U_leading_sign_16_0_rtn_not_nl));
  assign rtn = {IntLeadZero_16U_leading_sign_16_0_rtn_wrs_c_44_4_sdt_4 , (IntLeadZero_16U_leading_sign_16_0_rtn_IntLeadZero_16U_leading_sign_16_0_rtn_and_nl)};
  function [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input [0:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction
endmodule
//------> ./rtl.v
// ----------------------------------------------------------------------
// HLS HDL: Verilog Netlister
// HLS Version: 10.0/264918 Production Release
// HLS Date: Mon Aug 8 13:35:54 PDT 2016
//
// Generated by: ezhang@hk-sim-11-173
// Generated date: Mon Jun 12 22:24:10 2017
// ----------------------------------------------------------------------
//
// ------------------------------------------------------------------
// Design Unit: UINT16_TO_FP17_chn_o_rsci_unreg
// ------------------------------------------------------------------
module UINT16_TO_FP17_chn_o_rsci_unreg (
  in_0, outsig
);
  input in_0;
  output outsig;
// Interconnect Declarations for Component Instantiations
  assign outsig = in_0;
endmodule
// ------------------------------------------------------------------
// Design Unit: UINT16_TO_FP17_chn_a_rsci_unreg
// ------------------------------------------------------------------
module UINT16_TO_FP17_chn_a_rsci_unreg (
  in_0, outsig
);
  input in_0;
  output outsig;
// Interconnect Declarations for Component Instantiations
  assign outsig = in_0;
endmodule
// ------------------------------------------------------------------
// Design Unit: HLS_uint16_to_fp17_core_core_fsm
// FSM Module
// ------------------------------------------------------------------
module HLS_uint16_to_fp17_core_core_fsm (
  nvdla_core_clk, nvdla_core_rstn, core_wen, fsm_output
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input core_wen;
  output [1:0] fsm_output;
  reg [1:0] fsm_output;
// FSM State Type Declaration for HLS_uint16_to_fp17_core_core_fsm_1
  parameter
    core_rlp_C_0 = 1'd0,
    main_C_0 = 1'd1;
  reg [0:0] state_var;
  reg [0:0] state_var_NS;
// Interconnect Declarations for Component Instantiations
  always @(*)
  begin : HLS_uint16_to_fp17_core_core_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 2'b10;
        state_var_NS = main_C_0;
      end
// core_rlp_C_0
      default : begin
        fsm_output = 2'b1;
        state_var_NS = main_C_0;
      end
    endcase
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      state_var <= core_rlp_C_0;
    end
    else if ( core_wen ) begin
      state_var <= state_var_NS;
    end
  end
endmodule
// ------------------------------------------------------------------
// Design Unit: HLS_uint16_to_fp17_core_staller
// ------------------------------------------------------------------
module HLS_uint16_to_fp17_core_staller (
  nvdla_core_clk, nvdla_core_rstn, core_wen, chn_a_rsci_wen_comp, core_wten, chn_o_rsci_wen_comp
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output core_wen;
  input chn_a_rsci_wen_comp;
  output core_wten;
  reg core_wten;
  input chn_o_rsci_wen_comp;
// Interconnect Declarations for Component Instantiations
  assign core_wen = chn_a_rsci_wen_comp & chn_o_rsci_wen_comp;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      core_wten <= 1'b0;
    end
    else begin
      core_wten <= ~ core_wen;
    end
  end
endmodule
// ------------------------------------------------------------------
// Design Unit: HLS_uint16_to_fp17_core_chn_o_rsci_chn_o_wait_dp
// ------------------------------------------------------------------
module HLS_uint16_to_fp17_core_chn_o_rsci_chn_o_wait_dp (
  nvdla_core_clk, nvdla_core_rstn, chn_o_rsci_oswt, chn_o_rsci_bawt, chn_o_rsci_wen_comp,
      chn_o_rsci_biwt, chn_o_rsci_bdwt
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_o_rsci_oswt;
  output chn_o_rsci_bawt;
  output chn_o_rsci_wen_comp;
  input chn_o_rsci_biwt;
  input chn_o_rsci_bdwt;
// Interconnect Declarations
  reg chn_o_rsci_bcwt;
// Interconnect Declarations for Component Instantiations
  assign chn_o_rsci_bawt = chn_o_rsci_biwt | chn_o_rsci_bcwt;
  assign chn_o_rsci_wen_comp = (~ chn_o_rsci_oswt) | chn_o_rsci_bawt;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_o_rsci_bcwt <= 1'b0;
    end
    else begin
      chn_o_rsci_bcwt <= ~((~(chn_o_rsci_bcwt | chn_o_rsci_biwt)) | chn_o_rsci_bdwt);
    end
  end
endmodule
// ------------------------------------------------------------------
// Design Unit: HLS_uint16_to_fp17_core_chn_o_rsci_chn_o_wait_ctrl
// ------------------------------------------------------------------
module HLS_uint16_to_fp17_core_chn_o_rsci_chn_o_wait_ctrl (
  nvdla_core_clk, nvdla_core_rstn, chn_o_rsci_oswt, core_wen, core_wten, chn_o_rsci_iswt0,
      chn_o_rsci_ld_core_psct, chn_o_rsci_biwt, chn_o_rsci_bdwt, chn_o_rsci_ld_core_sct,
      chn_o_rsci_vd
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_o_rsci_oswt;
  input core_wen;
  input core_wten;
  input chn_o_rsci_iswt0;
  input chn_o_rsci_ld_core_psct;
  output chn_o_rsci_biwt;
  output chn_o_rsci_bdwt;
  output chn_o_rsci_ld_core_sct;
  input chn_o_rsci_vd;
// Interconnect Declarations
  wire chn_o_rsci_ogwt;
  wire chn_o_rsci_pdswt0;
  reg chn_o_rsci_icwt;
// Interconnect Declarations for Component Instantiations
  assign chn_o_rsci_pdswt0 = (~ core_wten) & chn_o_rsci_iswt0;
  assign chn_o_rsci_biwt = chn_o_rsci_ogwt & chn_o_rsci_vd;
  assign chn_o_rsci_ogwt = chn_o_rsci_pdswt0 | chn_o_rsci_icwt;
  assign chn_o_rsci_bdwt = chn_o_rsci_oswt & core_wen;
  assign chn_o_rsci_ld_core_sct = chn_o_rsci_ld_core_psct & chn_o_rsci_ogwt;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_o_rsci_icwt <= 1'b0;
    end
    else begin
      chn_o_rsci_icwt <= ~((~(chn_o_rsci_icwt | chn_o_rsci_pdswt0)) | chn_o_rsci_biwt);
    end
  end
endmodule
// ------------------------------------------------------------------
// Design Unit: HLS_uint16_to_fp17_core_chn_a_rsci_chn_a_wait_dp
// ------------------------------------------------------------------
module HLS_uint16_to_fp17_core_chn_a_rsci_chn_a_wait_dp (
  nvdla_core_clk, nvdla_core_rstn, chn_a_rsci_oswt, chn_a_rsci_bawt, chn_a_rsci_wen_comp,
      chn_a_rsci_d_mxwt, chn_a_rsci_biwt, chn_a_rsci_bdwt, chn_a_rsci_d
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_a_rsci_oswt;
  output chn_a_rsci_bawt;
  output chn_a_rsci_wen_comp;
  output [15:0] chn_a_rsci_d_mxwt;
  input chn_a_rsci_biwt;
  input chn_a_rsci_bdwt;
  input [15:0] chn_a_rsci_d;
// Interconnect Declarations
  reg chn_a_rsci_bcwt;
  reg [15:0] chn_a_rsci_d_bfwt;
// Interconnect Declarations for Component Instantiations
  assign chn_a_rsci_bawt = chn_a_rsci_biwt | chn_a_rsci_bcwt;
  assign chn_a_rsci_wen_comp = (~ chn_a_rsci_oswt) | chn_a_rsci_bawt;
  assign chn_a_rsci_d_mxwt = MUX_v_16_2_2(chn_a_rsci_d, chn_a_rsci_d_bfwt, chn_a_rsci_bcwt);
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_a_rsci_bcwt <= 1'b0;
      chn_a_rsci_d_bfwt <= 16'b0;
    end
    else begin
      chn_a_rsci_bcwt <= ~((~(chn_a_rsci_bcwt | chn_a_rsci_biwt)) | chn_a_rsci_bdwt);
      chn_a_rsci_d_bfwt <= chn_a_rsci_d_mxwt;
    end
  end
  function [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction
endmodule
// ------------------------------------------------------------------
// Design Unit: HLS_uint16_to_fp17_core_chn_a_rsci_chn_a_wait_ctrl
// ------------------------------------------------------------------
module HLS_uint16_to_fp17_core_chn_a_rsci_chn_a_wait_ctrl (
  nvdla_core_clk, nvdla_core_rstn, chn_a_rsci_oswt, core_wen, chn_a_rsci_iswt0, chn_a_rsci_ld_core_psct,
      core_wten, chn_a_rsci_biwt, chn_a_rsci_bdwt, chn_a_rsci_ld_core_sct, chn_a_rsci_vd
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_a_rsci_oswt;
  input core_wen;
  input chn_a_rsci_iswt0;
  input chn_a_rsci_ld_core_psct;
  input core_wten;
  output chn_a_rsci_biwt;
  output chn_a_rsci_bdwt;
  output chn_a_rsci_ld_core_sct;
  input chn_a_rsci_vd;
// Interconnect Declarations
  wire chn_a_rsci_ogwt;
  wire chn_a_rsci_pdswt0;
  reg chn_a_rsci_icwt;
// Interconnect Declarations for Component Instantiations
  assign chn_a_rsci_pdswt0 = (~ core_wten) & chn_a_rsci_iswt0;
  assign chn_a_rsci_biwt = chn_a_rsci_ogwt & chn_a_rsci_vd;
  assign chn_a_rsci_ogwt = chn_a_rsci_pdswt0 | chn_a_rsci_icwt;
  assign chn_a_rsci_bdwt = chn_a_rsci_oswt & core_wen;
  assign chn_a_rsci_ld_core_sct = chn_a_rsci_ld_core_psct & chn_a_rsci_ogwt;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_a_rsci_icwt <= 1'b0;
    end
    else begin
      chn_a_rsci_icwt <= ~((~(chn_a_rsci_icwt | chn_a_rsci_pdswt0)) | chn_a_rsci_biwt);
    end
  end
endmodule
// ------------------------------------------------------------------
// Design Unit: HLS_uint16_to_fp17_core_chn_o_rsci
// ------------------------------------------------------------------
module HLS_uint16_to_fp17_core_chn_o_rsci (
  nvdla_core_clk, nvdla_core_rstn, chn_o_rsc_z, chn_o_rsc_vz, chn_o_rsc_lz, chn_o_rsci_oswt,
      core_wen, core_wten, chn_o_rsci_iswt0, chn_o_rsci_bawt, chn_o_rsci_wen_comp,
      chn_o_rsci_ld_core_psct, chn_o_rsci_d
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output [16:0] chn_o_rsc_z;
  input chn_o_rsc_vz;
  output chn_o_rsc_lz;
  input chn_o_rsci_oswt;
  input core_wen;
  input core_wten;
  input chn_o_rsci_iswt0;
  output chn_o_rsci_bawt;
  output chn_o_rsci_wen_comp;
  input chn_o_rsci_ld_core_psct;
  input [16:0] chn_o_rsci_d;
// Interconnect Declarations
  wire chn_o_rsci_biwt;
  wire chn_o_rsci_bdwt;
  wire chn_o_rsci_ld_core_sct;
  wire chn_o_rsci_vd;
// Interconnect Declarations for Component Instantiations
  wire [16:0] nl_chn_o_rsci_d;
  assign nl_chn_o_rsci_d = {2'b0 , (chn_o_rsci_d[14:0])};
  UINT16_TO_FP17_mgc_out_stdreg_wait_v1 #(.rscid(32'sd2),
  .width(32'sd17)) chn_o_rsci (
      .ld(chn_o_rsci_ld_core_sct),
      .vd(chn_o_rsci_vd),
      .d(nl_chn_o_rsci_d[16:0]),
      .lz(chn_o_rsc_lz),
      .vz(chn_o_rsc_vz),
      .z(chn_o_rsc_z)
    );
  HLS_uint16_to_fp17_core_chn_o_rsci_chn_o_wait_ctrl HLS_uint16_to_fp17_core_chn_o_rsci_chn_o_wait_ctrl_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_o_rsci_oswt(chn_o_rsci_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .chn_o_rsci_iswt0(chn_o_rsci_iswt0),
      .chn_o_rsci_ld_core_psct(chn_o_rsci_ld_core_psct),
      .chn_o_rsci_biwt(chn_o_rsci_biwt),
      .chn_o_rsci_bdwt(chn_o_rsci_bdwt),
      .chn_o_rsci_ld_core_sct(chn_o_rsci_ld_core_sct),
      .chn_o_rsci_vd(chn_o_rsci_vd)
    );
  HLS_uint16_to_fp17_core_chn_o_rsci_chn_o_wait_dp HLS_uint16_to_fp17_core_chn_o_rsci_chn_o_wait_dp_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_o_rsci_oswt(chn_o_rsci_oswt),
      .chn_o_rsci_bawt(chn_o_rsci_bawt),
      .chn_o_rsci_wen_comp(chn_o_rsci_wen_comp),
      .chn_o_rsci_biwt(chn_o_rsci_biwt),
      .chn_o_rsci_bdwt(chn_o_rsci_bdwt)
    );
endmodule
// ------------------------------------------------------------------
// Design Unit: HLS_uint16_to_fp17_core_chn_a_rsci
// ------------------------------------------------------------------
module HLS_uint16_to_fp17_core_chn_a_rsci (
  nvdla_core_clk, nvdla_core_rstn, chn_a_rsc_z, chn_a_rsc_vz, chn_a_rsc_lz, chn_a_rsci_oswt,
      core_wen, chn_a_rsci_iswt0, chn_a_rsci_bawt, chn_a_rsci_wen_comp, chn_a_rsci_ld_core_psct,
      chn_a_rsci_d_mxwt, core_wten
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input [15:0] chn_a_rsc_z;
  input chn_a_rsc_vz;
  output chn_a_rsc_lz;
  input chn_a_rsci_oswt;
  input core_wen;
  input chn_a_rsci_iswt0;
  output chn_a_rsci_bawt;
  output chn_a_rsci_wen_comp;
  input chn_a_rsci_ld_core_psct;
  output [15:0] chn_a_rsci_d_mxwt;
  input core_wten;
// Interconnect Declarations
  wire chn_a_rsci_biwt;
  wire chn_a_rsci_bdwt;
  wire chn_a_rsci_ld_core_sct;
  wire chn_a_rsci_vd;
  wire [15:0] chn_a_rsci_d;
// Interconnect Declarations for Component Instantiations
  UINT16_TO_FP17_mgc_in_wire_wait_v1 #(.rscid(32'sd1),
  .width(32'sd16)) chn_a_rsci (
      .ld(chn_a_rsci_ld_core_sct),
      .vd(chn_a_rsci_vd),
      .d(chn_a_rsci_d),
      .lz(chn_a_rsc_lz),
      .vz(chn_a_rsc_vz),
      .z(chn_a_rsc_z)
    );
  HLS_uint16_to_fp17_core_chn_a_rsci_chn_a_wait_ctrl HLS_uint16_to_fp17_core_chn_a_rsci_chn_a_wait_ctrl_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_a_rsci_oswt(chn_a_rsci_oswt),
      .core_wen(core_wen),
      .chn_a_rsci_iswt0(chn_a_rsci_iswt0),
      .chn_a_rsci_ld_core_psct(chn_a_rsci_ld_core_psct),
      .core_wten(core_wten),
      .chn_a_rsci_biwt(chn_a_rsci_biwt),
      .chn_a_rsci_bdwt(chn_a_rsci_bdwt),
      .chn_a_rsci_ld_core_sct(chn_a_rsci_ld_core_sct),
      .chn_a_rsci_vd(chn_a_rsci_vd)
    );
  HLS_uint16_to_fp17_core_chn_a_rsci_chn_a_wait_dp HLS_uint16_to_fp17_core_chn_a_rsci_chn_a_wait_dp_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_a_rsci_oswt(chn_a_rsci_oswt),
      .chn_a_rsci_bawt(chn_a_rsci_bawt),
      .chn_a_rsci_wen_comp(chn_a_rsci_wen_comp),
      .chn_a_rsci_d_mxwt(chn_a_rsci_d_mxwt),
      .chn_a_rsci_biwt(chn_a_rsci_biwt),
      .chn_a_rsci_bdwt(chn_a_rsci_bdwt),
      .chn_a_rsci_d(chn_a_rsci_d)
    );
endmodule
// ------------------------------------------------------------------
// Design Unit: HLS_uint16_to_fp17_core
// ------------------------------------------------------------------
module HLS_uint16_to_fp17_core (
  nvdla_core_clk, nvdla_core_rstn, chn_a_rsc_z, chn_a_rsc_vz, chn_a_rsc_lz, chn_o_rsc_z,
      chn_o_rsc_vz, chn_o_rsc_lz, chn_a_rsci_oswt, chn_a_rsci_oswt_unreg, chn_o_rsci_oswt,
      chn_o_rsci_oswt_unreg
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input [15:0] chn_a_rsc_z;
  input chn_a_rsc_vz;
  output chn_a_rsc_lz;
  output [16:0] chn_o_rsc_z;
  input chn_o_rsc_vz;
  output chn_o_rsc_lz;
  input chn_a_rsci_oswt;
  output chn_a_rsci_oswt_unreg;
  input chn_o_rsci_oswt;
  output chn_o_rsci_oswt_unreg;
// Interconnect Declarations
  wire core_wen;
  reg chn_a_rsci_iswt0;
  wire chn_a_rsci_bawt;
  wire chn_a_rsci_wen_comp;
  reg chn_a_rsci_ld_core_psct;
  wire [15:0] chn_a_rsci_d_mxwt;
  wire core_wten;
  wire chn_o_rsci_bawt;
  wire chn_o_rsci_wen_comp;
  reg [4:0] chn_o_rsci_d_14_10;
  reg [9:0] chn_o_rsci_d_9_0;
  wire [1:0] fsm_output;
  wire and_dcpl_2;
  wire or_dcpl_1;
  wire and_dcpl_7;
  wire and_dcpl_22;
  wire or_tmp_7;
  reg FpMantRNE_17U_11U_else_and_svs;
  wire and_4_mdf;
  wire FpMantRNE_17U_11U_else_and_svs_mx1;
  wire FpFractionToFloat_16U_6U_10U_unequal_tmp;
  wire FpMantRNE_17U_11U_else_carry_sva;
  wire [16:0] FpMantRNE_17U_11U_i_data_sva;
  reg reg_chn_o_rsci_iswt0_cse;
  reg reg_chn_o_rsci_ld_core_psct_cse;
  wire or_cse;
  wire [10:0] FpMantRNE_17U_11U_else_ac_int_cctor_sva;
  wire [11:0] nl_FpMantRNE_17U_11U_else_ac_int_cctor_sva;
  wire nand_tmp;
  wire mux_tmp;
  wire chn_a_rsci_ld_core_psct_mx0c0;
  wire FpMantRNE_17U_11U_else_and_svs_mx0w0;
  wire FpFractionToFloat_16U_6U_10U_is_zero_lpi_1_dfm_1;
  wire [4:0] libraries_leading_sign_16_0_584ce9c19228fa5400845cefe3e6770649bb_1;
  wire FpFractionToFloat_16U_6U_10U_if_else_if_acc_itm_5_1;
  wire FpFractionToFloat_16U_6U_10U_if_else_else_if_acc_itm_4_1;
  wire[0:0] nor_9_nl;
  wire[0:0] nand_8_nl;
  wire[9:0] mux_4_nl;
  wire[0:0] and_53_nl;
  wire[4:0] and_nl;
  wire[4:0] mux_3_nl;
  wire[4:0] FpFractionToFloat_16U_6U_10U_nor_1_nl;
  wire[4:0] FpFractionToFloat_16U_6U_10U_if_else_else_else_acc_nl;
  wire[5:0] nl_FpFractionToFloat_16U_6U_10U_if_else_else_else_acc_nl;
  wire[0:0] FpFractionToFloat_16U_6U_10U_if_else_else_not_2_nl;
  wire[0:0] and_52_nl;
  wire[0:0] not_41_nl;
  wire[5:0] FpFractionToFloat_16U_6U_10U_if_else_if_acc_nl;
  wire[6:0] nl_FpFractionToFloat_16U_6U_10U_if_else_if_acc_nl;
  wire[4:0] FpFractionToFloat_16U_6U_10U_if_else_else_if_acc_nl;
  wire[5:0] nl_FpFractionToFloat_16U_6U_10U_if_else_else_if_acc_nl;
  wire[0:0] FpFractionToFloat_16U_6U_10U_if_else_mux_1_nl;
// Interconnect Declarations for Component Instantiations
  wire [6:0] nl_FpFractionToFloat_16U_6U_10U_if_shifted_frac_p1_lshift_rg_s;
  assign nl_FpFractionToFloat_16U_6U_10U_if_shifted_frac_p1_lshift_rg_s = conv_u2u_5_6(libraries_leading_sign_16_0_584ce9c19228fa5400845cefe3e6770649bb_1)
      + 6'b1;
  wire [16:0] nl_HLS_uint16_to_fp17_core_chn_o_rsci_inst_chn_o_rsci_d;
  assign nl_HLS_uint16_to_fp17_core_chn_o_rsci_inst_chn_o_rsci_d = {2'b0 , chn_o_rsci_d_14_10
      , chn_o_rsci_d_9_0};
  UINT16_TO_FP17_mgc_shift_l_v4 #(.width_a(32'sd16),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd17)) FpFractionToFloat_16U_6U_10U_if_shifted_frac_p1_lshift_rg (
      .a(chn_a_rsci_d_mxwt),
      .s(nl_FpFractionToFloat_16U_6U_10U_if_shifted_frac_p1_lshift_rg_s[5:0]),
      .z(FpMantRNE_17U_11U_i_data_sva)
    );
  UINT16_TO_FP17_leading_sign_16_0 leading_sign_16_0_rg (
      .mantissa(chn_a_rsci_d_mxwt),
      .rtn(libraries_leading_sign_16_0_584ce9c19228fa5400845cefe3e6770649bb_1)
    );
  HLS_uint16_to_fp17_core_chn_a_rsci HLS_uint16_to_fp17_core_chn_a_rsci_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_a_rsc_z(chn_a_rsc_z),
      .chn_a_rsc_vz(chn_a_rsc_vz),
      .chn_a_rsc_lz(chn_a_rsc_lz),
      .chn_a_rsci_oswt(chn_a_rsci_oswt),
      .core_wen(core_wen),
      .chn_a_rsci_iswt0(chn_a_rsci_iswt0),
      .chn_a_rsci_bawt(chn_a_rsci_bawt),
      .chn_a_rsci_wen_comp(chn_a_rsci_wen_comp),
      .chn_a_rsci_ld_core_psct(chn_a_rsci_ld_core_psct),
      .chn_a_rsci_d_mxwt(chn_a_rsci_d_mxwt),
      .core_wten(core_wten)
    );
  HLS_uint16_to_fp17_core_chn_o_rsci HLS_uint16_to_fp17_core_chn_o_rsci_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_o_rsc_z(chn_o_rsc_z),
      .chn_o_rsc_vz(chn_o_rsc_vz),
      .chn_o_rsc_lz(chn_o_rsc_lz),
      .chn_o_rsci_oswt(chn_o_rsci_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .chn_o_rsci_iswt0(reg_chn_o_rsci_iswt0_cse),
      .chn_o_rsci_bawt(chn_o_rsci_bawt),
      .chn_o_rsci_wen_comp(chn_o_rsci_wen_comp),
      .chn_o_rsci_ld_core_psct(reg_chn_o_rsci_ld_core_psct_cse),
      .chn_o_rsci_d(nl_HLS_uint16_to_fp17_core_chn_o_rsci_inst_chn_o_rsci_d[16:0])
    );
  HLS_uint16_to_fp17_core_staller HLS_uint16_to_fp17_core_staller_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .core_wen(core_wen),
      .chn_a_rsci_wen_comp(chn_a_rsci_wen_comp),
      .core_wten(core_wten),
      .chn_o_rsci_wen_comp(chn_o_rsci_wen_comp)
    );
  HLS_uint16_to_fp17_core_core_fsm HLS_uint16_to_fp17_core_core_fsm_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .core_wen(core_wen),
      .fsm_output(fsm_output)
    );
  assign nor_9_nl = ~(FpFractionToFloat_16U_6U_10U_if_else_if_acc_itm_5_1 | (~ FpMantRNE_17U_11U_else_and_svs_mx1));
  assign nand_8_nl = ~(FpFractionToFloat_16U_6U_10U_if_else_if_acc_itm_5_1 & FpMantRNE_17U_11U_else_and_svs_mx1);
  assign mux_tmp = MUX_s_1_2_2((nand_8_nl), (nor_9_nl), FpFractionToFloat_16U_6U_10U_if_else_else_if_acc_itm_4_1);
  assign nand_tmp = ~((~(FpMantRNE_17U_11U_else_and_svs_mx1 & (~ FpFractionToFloat_16U_6U_10U_if_else_if_acc_itm_5_1)))
      & FpFractionToFloat_16U_6U_10U_unequal_tmp);
  assign FpMantRNE_17U_11U_else_and_svs_mx0w0 = FpMantRNE_17U_11U_else_carry_sva
      & (FpMantRNE_17U_11U_i_data_sva[16:6]==11'b11111111111);
  assign FpMantRNE_17U_11U_else_and_svs_mx1 = MUX_s_1_2_2(FpMantRNE_17U_11U_else_and_svs_mx0w0,
      FpMantRNE_17U_11U_else_and_svs, and_dcpl_22);
  assign nl_FpFractionToFloat_16U_6U_10U_if_else_if_acc_nl = ({1'b1 , libraries_leading_sign_16_0_584ce9c19228fa5400845cefe3e6770649bb_1})
      + 6'b1;
  assign FpFractionToFloat_16U_6U_10U_if_else_if_acc_nl = nl_FpFractionToFloat_16U_6U_10U_if_else_if_acc_nl[5:0];
  assign FpFractionToFloat_16U_6U_10U_if_else_if_acc_itm_5_1 = readslicef_6_1_5((FpFractionToFloat_16U_6U_10U_if_else_if_acc_nl));
  assign nl_FpFractionToFloat_16U_6U_10U_if_else_else_if_acc_nl = ({1'b1 , (libraries_leading_sign_16_0_584ce9c19228fa5400845cefe3e6770649bb_1[4:1])})
      + 5'b1;
  assign FpFractionToFloat_16U_6U_10U_if_else_else_if_acc_nl = nl_FpFractionToFloat_16U_6U_10U_if_else_else_if_acc_nl[4:0];
  assign FpFractionToFloat_16U_6U_10U_if_else_else_if_acc_itm_4_1 = readslicef_5_1_4((FpFractionToFloat_16U_6U_10U_if_else_else_if_acc_nl));
  assign nl_FpMantRNE_17U_11U_else_ac_int_cctor_sva = (FpMantRNE_17U_11U_i_data_sva[16:6])
      + conv_u2u_1_11(FpMantRNE_17U_11U_else_carry_sva);
  assign FpMantRNE_17U_11U_else_ac_int_cctor_sva = nl_FpMantRNE_17U_11U_else_ac_int_cctor_sva[10:0];
  assign FpMantRNE_17U_11U_else_carry_sva = (FpMantRNE_17U_11U_i_data_sva[5]) & ((FpMantRNE_17U_11U_i_data_sva[0])
      | (FpMantRNE_17U_11U_i_data_sva[1]) | (FpMantRNE_17U_11U_i_data_sva[2]) | (FpMantRNE_17U_11U_i_data_sva[3])
      | (FpMantRNE_17U_11U_i_data_sva[4]) | (FpMantRNE_17U_11U_i_data_sva[6]));
  assign FpFractionToFloat_16U_6U_10U_unequal_tmp = (chn_a_rsci_d_mxwt!=16'b0000000000000000);
  assign FpFractionToFloat_16U_6U_10U_if_else_mux_1_nl = MUX_s_1_2_2(FpFractionToFloat_16U_6U_10U_if_else_else_if_acc_itm_4_1,
      FpFractionToFloat_16U_6U_10U_if_else_if_acc_itm_5_1, FpMantRNE_17U_11U_else_and_svs_mx1);
  assign FpFractionToFloat_16U_6U_10U_is_zero_lpi_1_dfm_1 = ~((FpFractionToFloat_16U_6U_10U_if_else_mux_1_nl)
      & FpFractionToFloat_16U_6U_10U_unequal_tmp);
  assign or_cse = chn_o_rsci_bawt | (~ reg_chn_o_rsci_ld_core_psct_cse);
  assign and_4_mdf = chn_a_rsci_bawt & or_cse;
  assign and_dcpl_2 = chn_o_rsci_bawt & reg_chn_o_rsci_ld_core_psct_cse;
  assign or_dcpl_1 = ~((~((~ chn_o_rsci_bawt) & reg_chn_o_rsci_ld_core_psct_cse))
      & chn_a_rsci_bawt);
  assign and_dcpl_7 = and_dcpl_2 & (~ chn_a_rsci_bawt);
  assign and_dcpl_22 = (chn_a_rsci_d_mxwt==16'b0000000000000000);
  assign or_tmp_7 = or_cse & chn_a_rsci_bawt & (fsm_output[1]);
  assign chn_a_rsci_ld_core_psct_mx0c0 = and_4_mdf | (fsm_output[0]);
  assign chn_a_rsci_oswt_unreg = or_tmp_7;
  assign chn_o_rsci_oswt_unreg = and_dcpl_2;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_a_rsci_iswt0 <= 1'b0;
      reg_chn_o_rsci_iswt0_cse <= 1'b0;
    end
    else if ( core_wen ) begin
      chn_a_rsci_iswt0 <= ~((~ and_4_mdf) & (fsm_output[1]));
      reg_chn_o_rsci_iswt0_cse <= or_tmp_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_a_rsci_ld_core_psct <= 1'b0;
    end
    else if ( core_wen & chn_a_rsci_ld_core_psct_mx0c0 ) begin
      chn_a_rsci_ld_core_psct <= chn_a_rsci_ld_core_psct_mx0c0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_o_rsci_d_9_0 <= 10'b0;
    end
    else if ( core_wen & (~(or_dcpl_1 | ((~(chn_o_rsci_bawt & reg_chn_o_rsci_ld_core_psct_cse
        & chn_a_rsci_bawt)) & (fsm_output[0])))) ) begin
      chn_o_rsci_d_9_0 <= (mux_4_nl) & (signext_10_1(~ mux_tmp)) & ({{9{FpFractionToFloat_16U_6U_10U_unequal_tmp}},
          FpFractionToFloat_16U_6U_10U_unequal_tmp}) & (signext_10_1(~ FpFractionToFloat_16U_6U_10U_is_zero_lpi_1_dfm_1));
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_o_rsci_d_14_10 <= 5'b0;
    end
    else if ( core_wen & (~(or_dcpl_1 | (fsm_output[0]))) ) begin
      chn_o_rsci_d_14_10 <= ~(MUX_v_5_2_2((and_nl), 5'b11111, FpFractionToFloat_16U_6U_10U_is_zero_lpi_1_dfm_1));
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_chn_o_rsci_ld_core_psct_cse <= 1'b0;
    end
    else if ( core_wen & (or_tmp_7 | and_dcpl_7) ) begin
      reg_chn_o_rsci_ld_core_psct_cse <= ~ and_dcpl_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMantRNE_17U_11U_else_and_svs <= 1'b0;
    end
    else if ( core_wen & (~(and_dcpl_22 | or_dcpl_1 | (fsm_output[0]))) ) begin
      FpMantRNE_17U_11U_else_and_svs <= FpMantRNE_17U_11U_else_and_svs_mx0w0;
    end
  end
  assign and_53_nl = FpMantRNE_17U_11U_else_and_svs_mx1 & (~ mux_tmp);
  assign mux_4_nl = MUX_v_10_2_2((FpMantRNE_17U_11U_else_ac_int_cctor_sva[9:0]),
      (FpMantRNE_17U_11U_else_ac_int_cctor_sva[10:1]), and_53_nl);
  assign nl_FpFractionToFloat_16U_6U_10U_if_else_else_else_acc_nl = (~ libraries_leading_sign_16_0_584ce9c19228fa5400845cefe3e6770649bb_1)
      + 5'b11111;
  assign FpFractionToFloat_16U_6U_10U_if_else_else_else_acc_nl = nl_FpFractionToFloat_16U_6U_10U_if_else_else_else_acc_nl[4:0];
  assign FpFractionToFloat_16U_6U_10U_if_else_else_not_2_nl = ~ FpFractionToFloat_16U_6U_10U_if_else_else_if_acc_itm_4_1;
  assign FpFractionToFloat_16U_6U_10U_nor_1_nl = ~(MUX_v_5_2_2((FpFractionToFloat_16U_6U_10U_if_else_else_else_acc_nl),
      5'b11111, (FpFractionToFloat_16U_6U_10U_if_else_else_not_2_nl)));
  assign and_52_nl = FpMantRNE_17U_11U_else_and_svs_mx1 & (~ nand_tmp);
  assign mux_3_nl = MUX_v_5_2_2((FpFractionToFloat_16U_6U_10U_nor_1_nl), libraries_leading_sign_16_0_584ce9c19228fa5400845cefe3e6770649bb_1,
      and_52_nl);
  assign not_41_nl = ~ nand_tmp;
  assign and_nl = MUX_v_5_2_2(5'b00000, (mux_3_nl), (not_41_nl));
  function [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction
  function [9:0] MUX_v_10_2_2;
    input [9:0] input_0;
    input [9:0] input_1;
    input [0:0] sel;
    reg [9:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_10_2_2 = result;
  end
  endfunction
  function [4:0] MUX_v_5_2_2;
    input [4:0] input_0;
    input [4:0] input_1;
    input [0:0] sel;
    reg [4:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_5_2_2 = result;
  end
  endfunction
  function [0:0] readslicef_5_1_4;
    input [4:0] vector;
    reg [4:0] tmp;
  begin
    tmp = vector >> 4;
    readslicef_5_1_4 = tmp[0:0];
  end
  endfunction
  function [0:0] readslicef_6_1_5;
    input [5:0] vector;
    reg [5:0] tmp;
  begin
    tmp = vector >> 5;
    readslicef_6_1_5 = tmp[0:0];
  end
  endfunction
  function [9:0] signext_10_1;
    input [0:0] vector;
  begin
    signext_10_1= {{9{vector[0]}}, vector};
  end
  endfunction
  function [10:0] conv_u2u_1_11 ;
    input [0:0] vector ;
  begin
    conv_u2u_1_11 = {{10{1'b0}}, vector};
  end
  endfunction
  function [5:0] conv_u2u_5_6 ;
    input [4:0] vector ;
  begin
    conv_u2u_5_6 = {1'b0, vector};
  end
  endfunction
endmodule
// ------------------------------------------------------------------
// Design Unit: HLS_uint16_to_fp17
// ------------------------------------------------------------------
module HLS_uint16_to_fp17 (
  nvdla_core_clk, nvdla_core_rstn, chn_a_rsc_z, chn_a_rsc_vz, chn_a_rsc_lz, chn_o_rsc_z,
      chn_o_rsc_vz, chn_o_rsc_lz
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input [15:0] chn_a_rsc_z;
  input chn_a_rsc_vz;
  output chn_a_rsc_lz;
  output [16:0] chn_o_rsc_z;
  input chn_o_rsc_vz;
  output chn_o_rsc_lz;
// Interconnect Declarations
  wire chn_a_rsci_oswt;
  wire chn_a_rsci_oswt_unreg;
  wire chn_o_rsci_oswt;
  wire chn_o_rsci_oswt_unreg;
// Interconnect Declarations for Component Instantiations
  UINT16_TO_FP17_chn_a_rsci_unreg chn_a_rsci_unreg_inst (
      .in_0(chn_a_rsci_oswt_unreg),
      .outsig(chn_a_rsci_oswt)
    );
  UINT16_TO_FP17_chn_o_rsci_unreg chn_o_rsci_unreg_inst (
      .in_0(chn_o_rsci_oswt_unreg),
      .outsig(chn_o_rsci_oswt)
    );
  HLS_uint16_to_fp17_core HLS_uint16_to_fp17_core_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_a_rsc_z(chn_a_rsc_z),
      .chn_a_rsc_vz(chn_a_rsc_vz),
      .chn_a_rsc_lz(chn_a_rsc_lz),
      .chn_o_rsc_z(chn_o_rsc_z),
      .chn_o_rsc_vz(chn_o_rsc_vz),
      .chn_o_rsc_lz(chn_o_rsc_lz),
      .chn_a_rsci_oswt(chn_a_rsci_oswt),
      .chn_a_rsci_oswt_unreg(chn_a_rsci_oswt_unreg),
      .chn_o_rsci_oswt(chn_o_rsci_oswt),
      .chn_o_rsci_oswt_unreg(chn_o_rsci_oswt_unreg)
    );
endmodule
